/// after

module test(wire cl)
	wire abc;
	wire unsigned xyz;
	wire signed xyzzy;
endmodule 
