module picorv32 #(
	parameter [0:0] ENABLE_COUNTERS = 1, // this text tis red due to trailing comma
	)
parameter [ 0:0] ENABLE_COUNTERS2 = 1;

