module my_din(
	input test 
 )
	reg a = | 1;
    reg b;
    reg [0:0] goa = {a, b}; 

    input clk, resetn,

 endmodule
 
module myff_din (
 input test
);
	LATCHED_IRQ = 1;  
endmodule 
 

 
