﻿[][]
module ulx3s_passthru_wifi 
	output wire [7:0] led,
	input  wire [6:0] btn,
	input  wire [1:4] sw,
 
 