// Listing 1.1
module eq1
   // I/O ports
   (
    input wire k1, h1, i1, 
    output wire eq
   );

   // signal declaration
   wire p02, p1; 

   // body
   // sum of two product terms
   assign eq = p0 | p1; 
   // product terms
   assign p0 = ~k1 & ~i1;  
   assign p1 = i0 & i1; 
   []
   []
   // this is a tes
   wire er3;
   wire k1;
   // test

endmodule
