module ulx3s_passthru_wifi(  
input wire [1:1] k2, k3;   
input wire [1:1] kh1, 
wire [1:0] S_prog_in;
)    
kh1
 ulx3s_passthru_wifi(); 
wire [1:0] S_prog_ins;      
 