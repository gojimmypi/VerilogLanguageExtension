module my_din (
    input [7:0] din
);

   din[7:0] == 0;
	din = 1;
endmodule  
  