module demo(
    inout v = 8 'h f_05, 
    inout a = 8'h f_05, 
    inout b = 8 'hf_05, 
    inout c = 8    'h  f_05, 
    inout bb = 3
)
v = 1;
endmodule
