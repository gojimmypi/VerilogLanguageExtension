// After

module other2(
  reg clk);

  wire a;
endmodule

module top(reg clk);
    other2 myOther(clk);
    myOther 
endmodule  




