
module picorv32 #(
	parameter [0:0] ENABLE_COUNTERS = 1,
	)
parameter [ 0:0] ENABLE_COUNTERS2 = 1;

